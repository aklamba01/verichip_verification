`timescale 1ns/1ps

`define SET_WRITE(addr,val,bytes)   \
   rw_ <= 1'b0;                     \
   chip_select <= 1'b1;             \
   byte_en <= bytes;                \
   address <= addr;                 \
   data_in <= val; 

`define SET_READ(addr)              \
   rw_ <= 1'b1;                     \
   chip_select <= 1'b1;             \
   byte_en <= 2'b00;                \
   address <= addr;                 \
   data_in <= 16'h0;

`define CLEAR_BUS                   \
   chip_select    <= 1'b0;          \
   address        <= 7'h0;          \
   byte_en        <= 2'h0;          \
   rw_            <= 1'b1;          \
   data_in        <= 16'h0; 

`define CLEAR_ALL                   \
   export_disable <= 1'b0;          \
   maroon         <= 1'b0;          \
   gold           <= 1'b0;          \
   `CLEAR_BUS

`define CHECK_VAL(val)              \
   if ( data_out != val )           \
       $display("bad read, got %h but expected %h at %t",data_out,val,$time());

`define CHECK_RW(addr,wval,rval,bytes)   \
  `WRITE_REG(addr,wval,bytes)            \
  `READ_REG(addr,rval)

`define CHIP_RESET                  \
   wait( clk == 1'b0 );             \	
   rst_b <= 1'b0;                   \
   wait( clk == 1'b1 );             \
   rst_b <= 1'b1;

// MR.C
`define READ_REG(addr,rval)	    \
   wait(clk == 1'b0);               \
   `SET_READ(addr)	               \
   wait(clk == 1'b1);               \
   `CHECK_VAL(rval)		            \
   `CLEAR_BUS                       \
   wait(clk == 1'b0);               

// MR.C
`define READ_REG_WITH_CS_OFF(addr, rval)  \
   wait(clk == 1'b0);                     \
   `SET_READ(addr)	                      \
   chip_select <= 1'b0;                   \
   wait(clk == 1'b1);                     \
   `CHECK_VAL(rval)		                    \
   `CLEAR_BUS                             \
   wait(clk == 1'b0);               

// MR.C
`define WRITE_REG(addr,wval,bytes)   \
   wait(clk == 1'b0);                \
   `SET_WRITE(addr,wval,bytes)       \
   wait(clk == 1'b1);                \
   `CLEAR_BUS                        \
   wait(clk == 1'b0);

// MR.C
`define WRITE_REG_WITH_CS_OFF(addr,wval,bytes)   \
   wait(clk == 1'b0);                \
   `SET_WRITE(addr,wval,bytes)       \
   chip_select <= 1'b0;              \
   wait(clk == 1'b1);                \
   `CLEAR_BUS                        \
   wait(clk == 1'b0);

// MR.C
`define TRANSITION_RST_TO_NORMAL    \
   `CLEAR_ALL                       \
   `CHIP_RESET                      \
   wait(clk == 1'b0);               \
   maroon <= 1'b0;                  \
   gold <= 1'b1;                    \
   wait(clk == 1'b1);               \
   `CLEAR_BUS                       \
   wait(clk == 1'b0);

// MR.C
`define ASSERT_MG                   \
   wait(clk == 1'b0);               \
   maroon <= 1'b1;                  \
   gold <= 1'b1;                    \
   wait(clk == 1'b1);               

// MR.C
`define ASSERT_M_NOT_G_NOT          \
   wait(clk == 1'b0);               \
   maroon <= 1'b0;                  \
   gold <= 1'b0;                    \
   wait(clk == 1'b1);               

// MR.C
`define ASSERT_M_G_NOT              \
   wait(clk == 1'b0);               \
   maroon <= 1'b1;                  \
   gold <= 1'b0;                    \
   wait(clk == 1'b1);               


// MR.C
`define TRANSITION_ERROR_TO_NORMAL    \
   wait(clk == 1'b0);               \
   maroon <= 1'b1;                  \
   gold <= 1'b0;                    \
   wait(clk == 1'b1);               \
   `CLEAR_BUS                       \
   wait(clk == 1'b0);

// MR.C
`define CHECK_STATE(state)          \
   `READ_CURRENT_STATE              \
   if(data_out[3:0] != state)       \
      $display("Current State: %h   \
      does NOT match the expected   \
      state: %h at %t!", data_out[3:0], state, $time());

// MR.C
`define READ_CURRENT_STATE          \
   `CLEAR_ALL                       \
   wait(clk == 1'b0);		            \
   `SET_READ(VCHIP_STA_ADDR)        \
   wait(clk == 1'b1);               \

// MR.C
`define TRANSITION_NORMAL_TO_ERROR                          \
   wait(clk == 1'b0);                                       \
   `SET_WRITE(VCHIP_CMD_ADDR, 16'h800F, BYTE_EN_MSB_LSB)    \
   wait(clk == 1'b1);                                       \    
   wait(clk == 1'b0);                                       \
   `SET_READ(VCHIP_STA_ADDR)                                \
   wait(clk == 1'b1);                    


// MR.C
//wait 1 cycle for operation TO BE WRITTEN TO CMD REGISTER
//wait 1 more cycle for OEPRATION TO EXECUTE
`define GENERATE_OVERFLOW                          \
   `CLEAR_ALL                                               \
   `WRITE_REG(VCHIP_ALU_LEFT_ADDR, 16'h7FFF, BYTE_EN_MSB_LSB)     \
   `WRITE_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001, BYTE_EN_MSB_LSB)     \
   wait(clk == 1'b0);                                       \
   `SET_WRITE(VCHIP_CMD_ADDR,VCHIP_ALU_VALID | VCHIP_ALU_ADD, BYTE_EN_MSB_LSB)    \
   wait(clk == 1'b1);                                       \    
   wait(clk == 1'b0);                                        \
   wait(clk == 1'b1);                                         \
   wait(clk == 1'b0);

//MR.C
`define EXECUTE_CMD(cmd, left_reg_val, right_reg_val)                      \
   //`CLEAR_ALL                                                              \
   `WRITE_REG(VCHIP_ALU_LEFT_ADDR, left_reg_val, BYTE_EN_MSB_LSB)          \
   `WRITE_REG(VCHIP_ALU_RIGHT_ADDR, right_reg_val, BYTE_EN_MSB_LSB)        \
   `WRITE_REG(VCHIP_CMD_ADDR,cmd, BYTE_EN_MSB_LSB)                         \
   wait(clk == 1'b1);                           


//MR.C
`define WAIT_CLK_CYCLE        \
   wait(clk == 1'b0);         \
   wait(clk == 1'b1);         

// RyUK
`define ASSERT_EXPORT_DISABLE       \
   export_disable <= 1'b1;

// RyUK
`define EXECUTE_BAD_COMMAND                                                        \
   `WRITE_REG(VCHIP_CMD_ADDR,VCHIP_ALU_MVL | VCHIP_ALU_VALID, BYTE_EN_MSB_LSB)     \

// RyUK
`define TRANSITION_NORMAL_TO_EXPORT       \
   wait(clk == 1'b0);		                  \
   `ASSERT_EXPORT_DISABLE                 \
   `EXECUTE_BAD_COMMAND                   \
   wait(clk == 1'b1);                     

  
    //Manz
`define TRANSITION_RST_TO_ERROR \
    `TRANSITION_RST_TO_NORMAL \
   `TRANSITION_NORMAL_TO_ERROR \
	
    
   
    

module top_verichip3 ();

logic clk;                       // system clock
logic rst_b;                     // chip reset
logic export_disable;            // disable features
logic interrupt_1;               // first interrupt
logic interrupt_2;               // second interrupt

logic maroon;                    // maroon state machine input
logic gold;                      // gold state machine input

logic chip_select;               // target of r/w
logic [6:0] address;             // address bus
logic [1:0] byte_en;             // write byte enables
logic       rw_;                 // read/write
logic [15:0] data_in;            // input data bus

logic [15:0] data_out;           // output data bus

logic [15:0] alu_left_random;
  logic [15:0] alu_right_random;
  logic [3:0] temp_state;
	
localparam VCHIP_VER_ADDR       = 7'h00;   // valid addresses
localparam VCHIP_STA_ADDR       = 7'h04;
localparam VCHIP_CMD_ADDR       = 7'h08;
localparam VCHIP_CON_ADDR       = 7'h0C;
localparam VCHIP_ALU_LEFT_ADDR  = 7'h10;
localparam VCHIP_ALU_RIGHT_ADDR = 7'h14;
localparam VCHIP_ALU_OUT_ADDR   = 7'h18;

localparam VCHIP_ALU_VALID = 16'h8000; // the valid bit
localparam VCHIP_ALU_ADD   = 16'h0001; // the various commands
localparam VCHIP_ALU_SUB   = 16'h0002; // OR the valid bit with the commands to do something
localparam VCHIP_ALU_MVL   = 16'h0003;
localparam VCHIP_ALU_MVR   = 16'h0004;
localparam VCHIP_ALU_SWA   = 16'h0005;
localparam VCHIP_ALU_SHL   = 16'h0006;
localparam VCHIP_ALU_SHR   = 16'h0007;

//RESET value for LEFT ALU REG
localparam VCHIP_ALU_LEFT_RST_VAL = 16'h0000;

//BYTE_EN 
localparam BYTE_EN_NONE = 2'b00;
localparam BYTE_EN_LSB = 2'b01;
localparam BYTE_EN_MSB = 2'b10;
localparam BYTE_EN_MSB_LSB = 2'b11;

//WRITE VALs to REGs
localparam ALL_ONE = 16'hFFFF;
localparam ALL_ZERO = 16'h0000;
localparam ALL_A = 16'hAAAA;
localparam ALL_5 = 16'h5555;

// States
localparam RESET_STATE = 4'h0;
localparam NORMAL_STATE = 4'h1;
localparam ERROR_STATE = 4'h2;
localparam EXPORT_VIOLATION_STATE = 4'h8;

// Undefined command
localparam UNDEFINED_CMD = 16'h000F;

initial      // get the clock running
begin
   clk <= 1'b0;
   while ( 1 )
   begin
      #5 clk <= 1'b1;
      #5 clk <= 1'b0;
   end
end

initial
begin
   // START WITH A NICE CLEAN INTERFACE AND A RESET
   `CLEAR_ALL
   `CHIP_RESET
   `CHECK_STATE(RESET_STATE)

// ADD TESTS HERE

///////NORMAL STATE////

//1 - ADD FUNCTIONALITY TEST IN NORMAL STATE -> 2 +ve no.
`TRANSITION_RST_TO_NORMAL
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h7FF0, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7FF0)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h7FF1)
`CHECK_STATE(NORMAL_STATE)


//2 - ADD OVERFLOW TEST IN NORMAL STATE -> +ve integers

`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h7FFF, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7FFF)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h8000)
`CHECK_STATE(ERROR_STATE)


//3 - ADD FUNCTIONALITY TEST IN NORMAL STATE -> a +ve and a -ve no.
`CLEAR_ALL
`CHIP_RESET
`TRANSITION_RST_TO_NORMAL
`WRITE_REG(VCHIP_ALU_OUT_ADDR, 16'h0001, BYTE_EN_MSB_LSB)          
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hFFF0, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hFFF0)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFF1)
`CHECK_STATE(NORMAL_STATE)

//4 - ADD OVERFLOW TEST IN NORMAL STATE -> -ve integers

`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h8000, 16'h8001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h8000)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h8001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0001)
`CHECK_STATE(ERROR_STATE)
  
  
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL 
`CHECK_STATE(NORMAL_STATE)
`ASSERT_EXPORT_DISABLE
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h7FFF, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7FFF)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h8000)
`CHECK_STATE(ERROR_STATE) 

///RESET STATE////

//5 - ADD FUNCTIONALITY TEST IN RESET STATE -> 2 +ve no.
`CLEAR_ALL
`CHIP_RESET
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h7FF0, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7FF0)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)

//6 - ADD OVERFLOW TEST IN RESET STATE -> +ve integers
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h7FFF, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7FFF)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)


//7 - ADD FUNCTIONALITY TEST IN RESET STATE -> a +ve and a -ve no.     
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hFFF0, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hFFF0)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)

//8 - ADD OVERFLOW TEST IN RESET STATE -> -ve integers
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h8000, 16'h8001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h8000)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h8001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)

//9. EXP Dis asserted, overflow
`ASSERT_EXPORT_DISABLE
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h7FFF, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7FFF)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)


///////////////////////////////// SUB FUNCTIONALITY TESTING /////////////////////////

/////////// SUB FUNCTIONALITY TESTING IN RESET STATE

// TEST: SUB +VE NUM FROM +VE NUM AND GENERATE +VE NUM
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h0003, 16'h0002)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0003)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0002) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)

// TEST: SUB A LARGE -VE NUMBER FROM +VE NUMBER: DOES NOT GENERATE OVERFLOW -> REMAINS IN RESET STATE
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h0001, 16'h8000)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0001)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h8000) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)


////////// SUB FUNCTIONALITY TESTING IN NORMAL STATE

// TEST: SUB 0 FROM +VE NUM
// SUB (5555) - (0) == (5555)
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h5555, 16'h0000)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h5555)
`CHECK_STATE(NORMAL_STATE)


// TEST: SUB +VE NUM FROM +VE NUM AND GENERATE +VE NUM
// SUB (+3) - (+2) == (1)
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h0003, 16'h0002)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0003)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0002) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0001)
`CHECK_STATE(NORMAL_STATE)

// TEST: SUB +VE NUM FROM +VE NUM AND GENERATE -VE NUM
// SUB (+2) - (+3) == (-1)
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h0002, 16'h0003)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0002)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0003) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
`CHECK_STATE(NORMAL_STATE)

// TEST: SUB A +VE NUMBER FROM -VE NUMBER TO GENERATE -VE NUM
// SUB (-1) - (+2) == (-3)
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'hFFFF, 16'h0002)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hFFFF)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0002) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFD)
`CHECK_STATE(NORMAL_STATE)

// TEST: SUB +VE NUM FROM -VE NUM GENERATING OVERFLOW -> MOVE TO ERROR STATE
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h8000, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h8000)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h7FFF)
`CHECK_STATE(ERROR_STATE)

// TEST: SUB A LARGE -VE NUMBER FROM +VE NUMBER TO GENERATE OVERFLOW -> MOVE TO ERROR STATE
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h0001, 16'h8000)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0001)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h8000) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h8001)
`CHECK_STATE(ERROR_STATE)

// TEST: SUB A SMALL -VE NUMBER FROM LARGE +VE NUMBER TO GENERATE OVERFLOW -> MOVE TO ERROR STATE
// SUB (7FFF) - (FFFF) == (8000)
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h7FFF, 16'hFFFF)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7FFF)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'hFFFF) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h8000)
`CHECK_STATE(ERROR_STATE)

// TEST: SUB A -VE NUMBER FROM +VE NUMBER TO GENERATE +VE NUM
// SUB (7000) - (FFFF) == (8001)
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h7000, 16'hFFFF)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7000)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'hFFFF) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h7001)
`CHECK_STATE(NORMAL_STATE)

// TEST: SUB A -VE NUMBER FROM -VE NUMBER TO GENERATE -VE NUM
// SUB (8000) - (FFFF) == (8001)
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h8000, 16'hFFFF)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h8000)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'hFFFF) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h8001)
`CHECK_STATE(NORMAL_STATE)

// TEST: SUB A -VE NUMBER FROM -VE NUMBER TO GENERATE +VE NUM
// SUB (FFFF) - (8000) == (7FFF)
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'hFFFF, 16'h8000)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hFFFF)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h8000) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h7FFF)
`CHECK_STATE(NORMAL_STATE)

/////////////////////////////////////////////////////////////////////////////////////

	
///////////////////////////////// SWAP FUNCTIONALITY TESTING ////////////////////////
// TEST 1: SWAP FUNCTIONALITY TESTS IN RESET STATE
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
//EXECUTE SWAP
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SWA, 16'hAAAA, 16'h5555)
//MAKE SURE THAT REGISTER VALUES ARE NOT SWAPPED
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)

// TEST 2: SWAP FUNCTIONALITY TESTS IN NORMAL STATE
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`CHECK_STATE(NORMAL_STATE)
//EXECUTE SWAP
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SWA, 16'hAAAA, 16'h5555)
//MAKE SURE THAT REGISTER VALUES ARE SWAPPED
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'hAAAA) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
`CHECK_STATE(NORMAL_STATE)
/////////////////////////////////////////////////////////////////////////////////////

  
/////////////////////////SHIFT FUNCTIONALITY TEST/////////////////////
///////////////////////// RESET -SHIFT LEFT //////////////////////////
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
  
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG - NEGATIVE
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - 0, Large Left 
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h5555, 16'h0000)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - < 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h5555, 16'h0006)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0006) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - > 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h5555, 16'h0016)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0016) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)


  
  
//EXECUTE SHIFT - 0, Small Left 
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h0005, 16'h0000)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0005)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - < 16, Small Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h0005, 16'h0004)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0005)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0004) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - > 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h0005, 16'h0014)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0005)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0014) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)  
  
//////////////////////////NORMAL - SHIFT LEFT///////////////////////// 
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
// TEST 2: SHIFT FUNCTIONALITY TESTS IN NORMAL STATE
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)

`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - 0, Large Left 
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h5555, 16'h0000)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000) 
//MAKE SURE THAT ALU_OUT IS THE SAME AS ALU LEFT
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h5555)
`CHECK_STATE(NORMAL_STATE)

  
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)   
//EXECUTE SHIFT - < 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h5555, 16'h0004)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0004) 
//MAKE SURE THAT ALU_OUT IS as expected
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h5550)
`CHECK_STATE(NORMAL_STATE)
  
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - > 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h5555, 16'h0016)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0016) 
//MAKE SURE THAT ALU_OUT IS as expected
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(NORMAL_STATE)


  
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - 0, Small Left 
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h0005, 16'h0000)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0005)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000) 
//MAKE SURE THAT ALU_OUT IS AS EXPECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0005)
`CHECK_STATE(NORMAL_STATE)

`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - < 16, Small Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h0005, 16'h0004)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0005)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0004) 
//MAKE SURE THAT ALU_OUT IS AS EXPECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0050)
`CHECK_STATE(NORMAL_STATE)

  
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - > 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h0005, 16'h0014)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0005)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0014) 
//MAKE SURE THAT ALU_OUT IS ALL ZERO 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(NORMAL_STATE) 

  
/////////////////////////SHIFT FUNCTIONALITY TEST/////////////////////
///////////////////////// RESET -SHIFT RIGHT //////////////////////////
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
  
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG - NEGATIVE
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - 0, Large Left 
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h5555, 16'h0000)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - < 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h5555, 16'h0006)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0006) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - > 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h5555, 16'h0016)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0016) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)


  
  
//EXECUTE SHIFT - 0, Small Left 
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h0005, 16'h0000)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0005)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - < 16, Small Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h0005, 16'h0004)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0005)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0004) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)
  
//EXECUTE SHIFT - > 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h0005, 16'h0014)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0005)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0014) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)  
  
//////////////////////////NORMAL - SHIFT RIGHT///////////////////////// 
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
// TEST 2: SHIFT FUNCTIONALITY TESTS IN NORMAL STATE
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)

`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - 0, Large Left 
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h5555, 16'h0000)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000) 
//MAKE SURE THAT ALU_OUT IS ALU LEFT
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h5555)
`CHECK_STATE(NORMAL_STATE)

  
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)   
//EXECUTE SHIFT - < 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h5555, 16'h0004)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0004) 
//MAKE SURE THAT ALU_OUT IS as expected
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0555)
`CHECK_STATE(NORMAL_STATE)
  
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - > 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h5555, 16'h0016)
//MAKE SURE THAT REGISTER VALUES ARE NT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0016) 
//MAKE SURE THAT ALU_OUT IS as expected
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(NORMAL_STATE)


  
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - 0, Small Left 
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h0050, 16'h0000)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0050)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000) 
//MAKE SURE THAT ALU_OUT IS ALU LEFT
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0050)
`CHECK_STATE(NORMAL_STATE)

`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - < 16, Small Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h0050, 16'h0004)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0050)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0004) 
//MAKE SURE THAT ALU_OUT IS AS EXPECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0005)
`CHECK_STATE(NORMAL_STATE)

  
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)  
//EXECUTE SHIFT - > 16, Small Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h0050, 16'h0014)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0050)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0014) 
//MAKE SURE THAT ALU_OUT IS ALL ZERO
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(NORMAL_STATE) 



///////////////////////////////// MOVE FUNCTIONALITY TESTING ////////////////////////
// TEST 1: MOVE FUNCTIONALITY TESTS IN RESET STATE
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)

//EXECUTE MOVE LEFT
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_MVL, 16'hAAAA, 16'h5555)
//MAKE SURE THAT LEFT & RIGHT REGISTERS ARE NOT AFFECTED
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)

//EXECUTE MOVE RIGHT
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_MVR, 16'hAAAA, 16'h5555)
//MAKE SURE THAT LEFT & RIGHT REGISTERS ARE NOT AFFECTED
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
`CHECK_STATE(RESET_STATE)


// TEST 2: MOVE FUNCTIONALITY TESTS IN NORMAL STATE
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`CHECK_STATE(NORMAL_STATE)

//EXECUTE MOVE LEFT
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_MVL, 16'hAAAA, 16'h5555)
//MAKE SURE THAT RIGHT REG IS NOT AFFECTED & LEFT CHANGES
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hFFFF)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
`CHECK_STATE(NORMAL_STATE)

//EXECUTE MOVE RIGHT
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_MVR, 16'hAAAA, 16'h5555)
//MAKE SURE THAT LEFT REG IS NOT AFFECTED & RIGHT CHANGES
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'hFFFF) 
//MAKE SURE THAT ALU_OUT IS NOT AFFECTED
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
`CHECK_STATE(NORMAL_STATE)

  for(int exp_dis = 0; exp_dis<2; exp_dis = exp_dis + 1)begin	
  	temp_state = RESET_STATE;
    	//$display("disable : %d", exp_dis);
  	for(logic [15:0] cmd = 16'h0000; cmd<=16'h800f; cmd = cmd + 1)begin
    	alu_left_random = $random();
  		alu_right_random = $random();
    	`CLEAR_ALL
		`CHIP_RESET
    	if(temp_state != RESET_STATE)begin
    		`TRANSITION_RST_TO_NORMAL
			`CHECK_STATE(NORMAL_STATE)
    	end
    	`CLEAR_BUS
      	`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555) 
    	if(temp_state != RESET_STATE)begin
      		`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
    	end
    	else begin 
      		`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
    	end
      	if (exp_dis == 1)begin
        	`ASSERT_EXPORT_DISABLE
      	end
        `CLEAR_BUS
    	`EXECUTE_CMD(cmd, alu_left_random, alu_right_random)
      	if (temp_state == EXPORT_VIOLATION_STATE)begin
          `READ_REG(VCHIP_ALU_LEFT_ADDR,16'h0000 )
          `READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000)
          `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
      	end
      	else begin 
			`READ_REG(VCHIP_ALU_LEFT_ADDR,alu_left_random )
			`READ_REG(VCHIP_ALU_RIGHT_ADDR, alu_right_random) 
        end 
      	if(temp_state ==  NORMAL_STATE || temp_state == ERROR_STATE)begin
      		`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
    	end
   		else begin 
          `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
    	end
   	`CHECK_STATE(temp_state)
	//$display(" %h, %d", cmd, temp_state);
    	if (cmd ==16'h000f)begin 
      		if(temp_state == RESET_STATE)begin
              cmd = 16'h7fff;
              //$display("Finished RESET invalid commands %d", exp_dis);
      		end
          	else begin
              cmd = 16'h8007;
              if(exp_dis == 1)begin 
                //$display("Started NORMAL invalid commands - EXP dis on");
              	temp_state = EXPORT_VIOLATION_STATE ;
              end
              else begin
                //$display("Started NORMAL invalid commands - EXP dis off");
                temp_state = ERROR_STATE;
              end 
      		end
    	end
      	if (cmd ==16'h800f)begin 
           if(temp_state == RESET_STATE)begin
             //$display("Finished RESET valid commands    %d", exp_dis);
              cmd = 16'hffff;
              temp_state = NORMAL_STATE;
           end
        end
  	end
  end
  //NO OP WITH EXP DISABLE WITH AND WITHOUT VALID
 `CLEAR_ALL
 `CHIP_RESET
 `TRANSITION_RST_TO_NORMAL
  alu_left_random = $random();
  alu_right_random = $random();
  `EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555) 
 `READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
 `ASSERT_EXPORT_DISABLE
 `EXECUTE_CMD(16'h8000, alu_left_random, alu_right_random)
 `READ_REG(VCHIP_ALU_LEFT_ADDR, alu_left_random)
 `READ_REG(VCHIP_ALU_RIGHT_ADDR, alu_right_random)
 `READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
 `CHECK_STATE(NORMAL_STATE)


 `CLEAR_ALL
 `CHIP_RESET
 `TRANSITION_RST_TO_NORMAL
  alu_left_random = $random();
  alu_right_random = $random();
  `EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5554) 
 `READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFE)
 `ASSERT_EXPORT_DISABLE
 `EXECUTE_CMD(16'h0000, alu_left_random, alu_right_random)
 `READ_REG(VCHIP_ALU_LEFT_ADDR, alu_left_random)
 `READ_REG(VCHIP_ALU_RIGHT_ADDR, alu_right_random)
 `READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFE)
 `CHECK_STATE(NORMAL_STATE)

//

//NO OP WITHOUT EXP DISABLE WITH AND WITHOUT VALID
 `CLEAR_ALL
 `CHIP_RESET
 `TRANSITION_RST_TO_NORMAL
  alu_left_random = $random();
  alu_right_random = $random();
  `EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555) 
 `READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
 `EXECUTE_CMD(16'h8000, alu_left_random, alu_right_random)
 `READ_REG(VCHIP_ALU_LEFT_ADDR, alu_left_random)
 `READ_REG(VCHIP_ALU_RIGHT_ADDR, alu_right_random)
 `READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
 `CHECK_STATE(NORMAL_STATE)


 `CLEAR_ALL
 `CHIP_RESET
 `TRANSITION_RST_TO_NORMAL
  alu_left_random = $random();
  alu_right_random = $random();
  `EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5554) 
 `READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFE)
 
 `EXECUTE_CMD(16'h0000, alu_left_random, alu_right_random)
 `READ_REG(VCHIP_ALU_LEFT_ADDR, alu_left_random)
 `READ_REG(VCHIP_ALU_RIGHT_ADDR, alu_right_random)
 `READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFE)
 `CHECK_STATE(NORMAL_STATE)

//
//7. NORMAL STATE - SHIFT LEFT by 11 bits
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)   
//EXECUTE SHIFT - < 16, Large Left
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHL, 16'h5555, 16'h000b)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h000b) 
//MAKE SURE THAT ALU_OUT IS as expected
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'ha800)
`CHECK_STATE(NORMAL_STATE)


// ADD TO CHECK CARRY 
`CLEAR_ALL
`CHIP_RESET
`TRANSITION_RST_TO_NORMAL
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h3fff, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h3fff)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h4000)
`CHECK_STATE(NORMAL_STATE)

//ADD 2 -ve NUMBERS
`CLEAR_ALL
`CHIP_RESET
`TRANSITION_RST_TO_NORMAL
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hff88, 16'hffff)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hff88)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'hffff) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hff87)
`CHECK_STATE(NORMAL_STATE)

//Subtract to generate overflow with export_disable asserted!
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`ASSERT_EXPORT_DISABLE
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h8000, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h8000)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h7FFF)
`CHECK_STATE(ERROR_STATE)

//Subtract with BORROW case
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
//EXECUTE ADD CMD TO WRITE NON-ZERO VALUE TO ALU OUT REG
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h7000, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7000)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h6FFF)
`CHECK_STATE(NORMAL_STATE)


//COMMANDS 3-F FOR EXPORT DISABLE ASSERTED 
for (logic[15:0] cmd = 16'h0003; cmd <= 16'h000F; cmd = cmd + 1 )
begin
   `ASSERT_EXPORT_DISABLE
   `EXECUTE_CMD(VCHIP_ALU_VALID | cmd, 16'hAAAA, 16'h5555)
   //CHECK REG VALS
   `READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0000)
   `READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0000)
   `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)
   `CHECK_STATE(EXPORT_VIOLATION_STATE)
   `CHIP_RESET
   `CHECK_STATE(RESET_STATE)
   `TRANSITION_RST_TO_NORMAL
   `CHECK_STATE(NORMAL_STATE)
end

//COMMAND 1 and 2 WITH EXPORT DISABLE ASSERTED

//ADD FUNCTIONALITY TEST IN NORMAL STATE with EXPORT -> 2 +ve no.
`CHIP_RESET
`TRANSITION_RST_TO_NORMAL
`ASSERT_EXPORT_DISABLE
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'h7FF0, 16'h0001)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h7FF0)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0001) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h7FF1)
`CHECK_STATE(NORMAL_STATE)

// TEST: SUB +VE NUM FROM +VE NUM AND GENERATE +VE NUM
// SUB (+3) - (+2) == (1)
`CLEAR_ALL
`CHIP_RESET
`CHECK_STATE(RESET_STATE)
`TRANSITION_RST_TO_NORMAL
`CHECK_STATE(NORMAL_STATE)
`ASSERT_EXPORT_DISABLE
//EXECUTE SUB
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SUB, 16'h0003, 16'h0002)
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h0003)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h0002) 
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0001)
`CHECK_STATE(NORMAL_STATE)

  
//7. NORMAL STATE - SHIFT RIGHT by 11 bits
`EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_ADD, 16'hAAAA, 16'h5555)
`READ_REG(VCHIP_ALU_OUT_ADDR, 16'hFFFF)   
//EXECUTE SHIFT - < 16, Large Left
  `EXECUTE_CMD(VCHIP_ALU_VALID | VCHIP_ALU_SHR, 16'h5555, 16'h000b)
//MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
`READ_REG(VCHIP_ALU_LEFT_ADDR, 16'h5555)
`READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h000b) 
//MAKE SURE THAT ALU_OUT IS as expected
  `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h000a)
`CHECK_STATE(NORMAL_STATE)

//////NORMAL STATE LOOPS////
///////// valid bit missing //////
for(logic[15:0] cmd = 16'h0000; cmd <= 16'h000F; cmd = cmd +1)
begin
    `CHECK_STATE(NORMAL_STATE)
    `EXECUTE_CMD(cmd, 16'hAAAA, 16'h5555)
    //MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
    `READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
    `READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
    `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h000a)  
    `CHECK_STATE(NORMAL_STATE)
end

///////// valid bit missing //////
for(logic[15:0] cmd = 16'h0000; cmd <= 16'h000F; cmd = cmd +1)
begin
    `CHECK_STATE(NORMAL_STATE)
    `ASSERT_EXPORT_DISABLE
    `EXECUTE_CMD(cmd, 16'hAAAA, 16'h5555)
    //MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
    `READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
    `READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
    `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h000a)  
    `CHECK_STATE(NORMAL_STATE)
end



/////END OF NORMAL STATE LOOPS////


////////RESET STATE LOOPS///////
`CLEAR_ALL
`CHIP_RESET
///////// valid bit missing in reset //////
for(logic[15:0] cmd = 16'h0000; cmd <= 16'h000F; cmd = cmd +1)
begin
   
    `CHECK_STATE(RESET_STATE)
    `EXECUTE_CMD(cmd, 16'hAAAA, 16'h5555)
    //MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
    `READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
    `READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
    `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)  
    `CHECK_STATE(RESET_STATE)
end

///////// valid bit not missing in reset //////
for(logic[15:0] cmd = 16'h8000; cmd <= 16'h800f; cmd = cmd +1)
begin
   
    `CHECK_STATE(RESET_STATE)
    `EXECUTE_CMD(cmd, 16'hAAAA, 16'h5555)
    //MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
    `READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
    `READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
    `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)  
    `CHECK_STATE(RESET_STATE)
end

///////// valid bit missing in reset - expo disable //////
for(logic[15:0] cmd = 16'h0000; cmd <= 16'h000F; cmd = cmd +1)
begin
   
    `CHECK_STATE(RESET_STATE)
    `ASSERT_EXPORT_DISABLE
    `EXECUTE_CMD(cmd, 16'hAAAA, 16'h5555)
    //MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
    `READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
    `READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
    `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)  
    `CHECK_STATE(RESET_STATE)
end

///////// valid bit not missing in reset - expo disable//////
for(logic[15:0] cmd = 16'h8000; cmd <= 16'h800f; cmd = cmd +1)
begin
   
    `CHECK_STATE(RESET_STATE)
    `ASSERT_EXPORT_DISABLE
    `EXECUTE_CMD(cmd, 16'hAAAA, 16'h5555)
    //MAKE SURE THAT REGISTER VALUES ARE NOT ALTERED 
    `READ_REG(VCHIP_ALU_LEFT_ADDR, 16'hAAAA)
    `READ_REG(VCHIP_ALU_RIGHT_ADDR, 16'h5555) 
    `READ_REG(VCHIP_ALU_OUT_ADDR, 16'h0000)  
    `CHECK_STATE(RESET_STATE)
end


// MUST LEAVE SO GRADING WORKS!
   wait(clk == 1'b0);   
   wait(clk == 1'b1);
   wait(clk == 1'b0);
   $finish; // THIS MUST BE THE LAST THING YOU EXECUTE!
end // initial begin

// instantiate the VeriChip!
verichip3 verichip3 (.clk           ( clk            ),    // system clock
                   .rst_b         ( rst_b          ),    // chip reset
                   .export_disable( export_disable ),    // disable features
                   .interrupt_1   ( interrupt_1    ),    // first interrupt
                   .interrupt_2   ( interrupt_2    ),    // second interrupt
 
                   .maroon        ( maroon         ),    // maroon state machine input
                   .gold          ( gold           ),    // gold state machine input

                   .chip_select   ( chip_select    ),    // target of r/w
                   .address       ( address        ),    // address bus
                   .byte_en       ( byte_en        ),    // write byte enables
                   .rw_           ( rw_            ),    // read/write
                   .data_in       ( data_in        ),    // data bus

                   .data_out      ( data_out       ) );  // output data bus

endmodule // top_verichip
